library verilog;
use verilog.vl_types.all;
entity g21_7_segment_decoder_vlg_vec_tst is
end g21_7_segment_decoder_vlg_vec_tst;
