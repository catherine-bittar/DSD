library verilog;
use verilog.vl_types.all;
entity g21_lab2_vlg_vec_tst is
end g21_lab2_vlg_vec_tst;
