library verilog;
use verilog.vl_types.all;
entity g21_dealer_FSM_vlg_vec_tst is
end g21_dealer_FSM_vlg_vec_tst;
