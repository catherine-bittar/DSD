library verilog;
use verilog.vl_types.all;
entity g21_SPG_vlg_vec_tst is
end g21_SPG_vlg_vec_tst;
