library verilog;
use verilog.vl_types.all;
entity g21_test_bed_lab4_vlg_vec_tst is
end g21_test_bed_lab4_vlg_vec_tst;
