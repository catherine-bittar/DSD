library verilog;
use verilog.vl_types.all;
entity g21_pop_enable_vlg_vec_tst is
end g21_pop_enable_vlg_vec_tst;
