library verilog;
use verilog.vl_types.all;
entity g21_dealer_FSM_vlg_check_tst is
    port(
        Rand_Enable     : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g21_dealer_FSM_vlg_check_tst;
